interface spi_if;
    logic i_sclk;
    logic spi_cs_n;
    logic spi_mosi;
    logic spi_miso;
endinterface
