/**
 * SPI to AXI Stream Bridge
 * 
 * Simple bridge that streams SPI data directly to AXI Stream interface
 * Uses IMPLICIT_FRAMING mode - axis_wb_master detects command bytes (0xA1/0xA2)
 * 
 * Operation:
 * 1. SPI bytes are forwarded directly to AXI Stream
 * 2. axis_wb_master looks for READ_REQ (0xA1) or WRITE_REQ (0xA2) to detect frame start
 * 3. Command format defines packet length, so tlast is not needed
 * 4. Responses are streamed back to SPI
 */

module spi_axis_adapter #(
    parameter AXIS_DATA_WIDTH = 8
) (
    input  logic                       clk,
    input  logic                       rst_n,
    
    // SPI Slave Interface
    input  logic [7:0]                 spi_rx_data,
    input  logic                       spi_rx_valid,
    output logic [7:0]                 spi_tx_data,
    output logic                       spi_tx_valid,
    input  logic                       spi_busy,
    input  logic                       spi_cs_n,      // Optional: can be used for debug/status
    
    // AXI Stream Output (to axis_wb_master input)
    output logic [AXIS_DATA_WIDTH-1:0] m_axis_tdata,
    output logic                       m_axis_tvalid,
    input  logic                       m_axis_tready,
    output logic                       m_axis_tlast,  // Not used in implicit framing
    
    // AXI Stream Input (from axis_wb_master output)
    input  logic [AXIS_DATA_WIDTH-1:0] s_axis_tdata,
    input  logic                       s_axis_tvalid,
    output logic                       s_axis_tready,
    input  logic                       s_axis_tlast
);

    // =============================
    // SPI RX to AXI Stream TX
    // Simple pass-through
    // =============================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            m_axis_tdata <= 8'h0;
            m_axis_tvalid <= 1'b0;
        end else begin
            // Clear valid when data is accepted
            if (m_axis_tvalid && m_axis_tready) begin
                m_axis_tvalid <= 1'b0;
            end
            
            // Forward SPI RX data to AXI Stream
            if (spi_rx_valid && !m_axis_tvalid) begin
                m_axis_tdata <= spi_rx_data;
                m_axis_tvalid <= 1'b1;
            end
        end
    end
    
    // tlast not used in implicit framing mode
    assign m_axis_tlast = 1'b0;
    
    // =============================
    // AXI Stream RX to SPI TX
    // Simple pass-through
    // =============================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            spi_tx_data <= 8'h0;
            spi_tx_valid <= 1'b0;
            s_axis_tready <= 1'b1;
        end else begin
            spi_tx_valid <= 1'b0;
            s_axis_tready <= 1'b1;  // Always ready to receive
            
            // Forward AXI Stream data to SPI TX when not busy
            if (s_axis_tvalid && s_axis_tready && !spi_busy) begin
                spi_tx_data <= s_axis_tdata;
                spi_tx_valid <= 1'b1;
            end
        end
    end

endmodule
    
    // =============================
    // AXI Stream RX to SPI TX
    // =============================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            spi_tx_data <= 8'h0;
            spi_tx_valid <= 1'b0;
            s_axis_tready <= 1'b1;  // Always ready to receive
        end else begin
            spi_tx_valid <= 1'b0;
            s_axis_tready <= 1'b1;
            
            // Forward AXI Stream data to SPI TX
            if (s_axis_tvalid && s_axis_tready && !spi_busy) begin
                spi_tx_data <= s_axis_tdata;
                spi_tx_valid <= 1'b1;
            end
        end
    end

endmodule
