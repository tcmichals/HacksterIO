module spi_slave #(
    parameter DATA_WIDTH = 8
)(
    input  logic                   i_clk,
    input  logic                   i_rst,
    
    // SPI Physical Interface
    input  logic                   i_sclk,
    input  logic                   i_cs_n,
    input  logic                   i_mosi,
    output logic                   o_miso,
    
    // User / System Interface
    input  logic [DATA_WIDTH-1:0]  i_tx_data,  // Data to send
    input  logic                   i_tx_valid, // Pulse high to load data
    output logic                   o_tx_ready, // High = Safe to load new data
    output logic                   o_busy,     // High = SPI transaction in progress
    
    output logic [DATA_WIDTH-1:0]  o_rx_data,  // Received data
    output logic                   o_data_valid // High = New rx_data available
);

    // --- 1. Synchronization & Edge Detection ---
    logic [2:0] sclk_sync;
    logic [2:0] cs_n_sync;
    logic [1:0] mosi_sync;

    always_ff @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            sclk_sync <= 3'b000;
            cs_n_sync <= 3'b111;
            mosi_sync <= 2'b00;
        end else begin
            sclk_sync <= {sclk_sync[1:0], i_sclk};
            cs_n_sync <= {cs_n_sync[1:0], i_cs_n};
            mosi_sync <= {mosi_sync[0], i_mosi};
        end
    end

    // Derived signals from synchronizers
    wire sclk_rising  = (sclk_sync[2:1] == 2'b01);
    wire sclk_falling = (sclk_sync[2:1] == 2'b10);
    wire cs_active    = ~cs_n_sync[1]; // Active Low CS
    
    // Output the Busy status immediately based on synchronized CS
    assign o_busy = cs_active;

    // --- 2. Data Path & Logic ---
    logic [$clog2(DATA_WIDTH)-1:0] bit_cnt;
    logic [DATA_WIDTH-1:0] rx_shift_reg;
    logic [DATA_WIDTH-1:0] tx_shift_reg;
    logic [DATA_WIDTH-1:0] tx_holding_reg; 

    always_ff @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            bit_cnt        <= DATA_WIDTH - 1;
            o_rx_data      <= '0;
            o_data_valid   <= 1'b0;
            rx_shift_reg   <= '0;
            tx_shift_reg   <= '0;
            tx_holding_reg <= '0;
            o_tx_ready     <= 1'b1;
        end else begin
            o_data_valid <= 1'b0;

            // --- A. User Interface Logic (Safe Loading) ---
            if (i_tx_valid && o_tx_ready) begin
                tx_holding_reg <= i_tx_data;
                o_tx_ready     <= 1'b0; // Lock buffer until SPI takes it
            end

            // --- B. SPI Transaction Logic ---
            if (!cs_active) begin
                // IDLE STATE
                bit_cnt <= DATA_WIDTH - 1; 
                
                // If the user loaded data, move it to the shifter immediately
                if (o_tx_ready == 1'b0) begin
                    tx_shift_reg <= tx_holding_reg;
                    o_tx_ready   <= 1'b1; // Unlock buffer
                end
            end 
            else begin
                // ACTIVE STATE (Busy)
                
                // Sample MOSI (Rising Edge)
                if (sclk_rising) begin
                    rx_shift_reg <= {rx_shift_reg[DATA_WIDTH-2:0], mosi_sync[1]};
                    if (bit_cnt == 0) begin
                        o_rx_data    <= {rx_shift_reg[DATA_WIDTH-2:0], mosi_sync[1]};
                        o_data_valid <= 1'b1;
                    end
                end

                // Shift MISO (Falling Edge)
                if (sclk_falling) begin
                    if (bit_cnt > 0) begin
                        bit_cnt      <= bit_cnt - 1;
                        tx_shift_reg <= {tx_shift_reg[DATA_WIDTH-2:0], 1'b0};
                    end else begin
                        // Byte complete. Prepare for next byte in stream (if any).
                        bit_cnt <= DATA_WIDTH - 1;
                        
                        // Check if user provided new data in holding register
                        if (o_tx_ready == 1'b0) begin
                            tx_shift_reg <= tx_holding_reg;
                            o_tx_ready   <= 1'b1; // Unlock buffer
                        end else begin
                            tx_shift_reg <= '0; // Underflow: Send Zeros
                        end
                    end
                end
            end
        end
    end

    // Tri-state MISO
    assign o_miso = (cs_active) ? tx_shift_reg[DATA_WIDTH-1] : 1'bZ;

endmodule // SPI_Slave